package AHB5_Slave_package;
  `include "../sv/AHB5_Slave_Transaction.sv"
  `include "../sv/AHB5_Slave_Configuration.sv"
  `include "../sv/AHB5_Slave_generator.sv"
  `include "../sv/AHB5_Slave_Driver.sv"
  `include "../sv/AHB5_Slave_Monitor.sv"
  `include "../sv/AHB5_Slave_Scoreboard.sv"
  `include "../sve/AHB5_Slave_Dummy_master.sv"

endpackage


`include "../sv/AHB5_Slave_interface.sv"
