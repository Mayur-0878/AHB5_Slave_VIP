class configure;
 parameter size=8;
 
 bit mem[];
 


endclass
