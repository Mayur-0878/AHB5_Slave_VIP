package AHB5_Slave_package;
  `include "../sv/AHB5_Slave_Transaction.sv"
  `include "../sv/AHB5_Slave_generator.sv"
  `include "../sv/AHB5_Slave_Driver.sv"
  `include "../sv/AHB5_Slave_Monitor.sv"
  `include "../sv/AHB5_Slave_Scoreboard.sv"
  `include "../sv/AHB5_Slave_Dummy_master.sv"
  `include "../sv/AHB5_Slave_Environment.sv"
  `include "../sve/AHB5_Slave_Configuration.sv"
  `include "../sve/AHB5_Slave_test.sv"
  `include "AHB5_Slave_top.sv"


endpackage
